module Main(
	CLK50,
	PAUSE_KEY,
	STOP_KEY,
	RATIO_SW,
	RECORD_SW,
	NORMAL_SPEED_SW,
);
	Clock c1();
endmodule
